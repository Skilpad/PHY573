
library IEEE;
use IEEE.std_logic_1164.all;

entity afficheur_hexa is
port(

-- A faire

);
end afficheur_hexa;


architecture afficheur_hexa_arch of afficheur_hexa is
begin

-- A faire

end afficheur_hexa_arch;