
library IEEE;
use IEEE.std_logic_1164.all;

entity generateur_coefs is
port(

-- A faire

);
end generateur_coefs;


architecture generateur_coefs_arch of generateur_coefs is
begin

-- A faire

end generateur_coefs_arch;